LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ssegNEW IS
	PORT( bcd	: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
			neg 	: IN STD_LOGIC;
			leds 	: OUT STD_LOGIC_VECTOR(1 TO 7);
			ledss : OUT STD_LOGIC_VECTOR(1 TO 7));
END ssegNEW;
			
ARCHITECTURE Behavior OF ssegNEW IS
BEGIN
	PROCESS(bcd)
	BEGIN	
		CASE bcd IS					-- abcdefg
			WHEN "0000" => leds <= "1111110";
			WHEN "0001" => leds <= "0110000"; --y
			WHEN "0010" => leds <= "1101101";
			WHEN "0011" => leds <= "1111001";--y
			WHEN "0100" => leds <= "0110011";
			WHEN "0101" => leds <= "1011011";--y
			WHEN "0110" => leds <= "1011111";
			WHEN "0111" => leds <= "1110000";--y
			WHEN "1000" => leds <= "1111111";
			WHEN "1001" => leds <= "1110011";--y
			WHEN "1010" => leds <= "1110111"; --A 
			WHEN "1011" => leds <= "0011111"; --B(y)
			WHEN "1100" => leds <= "1001110"; --C
			WHEN "1101" => leds <= "0111101"; --D(y)
			WHEN "1110" => leds <= "1001111"; --E
			WHEN "1111" => leds <= "1000111"; --F(y)
			WHEN OTHERS => leds <= "-------";
		END CASE;
	END PROCESS;
	
	PROCESS (neg)
	BEGIN
		IF(neg = '1') THEN
		ledss <= "0000001";
		
		ELSE
		ledss <= "0000000";
	END IF;
	END PROCESS;
END Behavior;
